library verilog;
use verilog.vl_types.all;
entity Register_file_tb is
end Register_file_tb;
